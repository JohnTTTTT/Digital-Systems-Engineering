module Datapath (input clk, CU_clk, Reset, Stop,
					  output [31:0] Busout);
	endmodule
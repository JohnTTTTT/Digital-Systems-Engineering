module ROR (input [31:0] a, b, output[31:0] result);
	reg [31:0] res;
	assign result = res;
	always @(a or b) begin
		case (b)
				5'd1:	res <= {a[0], a[31:1]};
				5'd2:	res <= {a[1:0], a[31:2]};
				5'd3:	res <= {a[2:0], a[31:3]};
				5'd4:	res <= {a[3:0], a[31:4]};
				5'd5:	res <= {a[4:0], a[31:5]};
				5'd6:	res <= {a[5:0], a[31:6]};
				5'd7:	res <= {a[6:0], a[31:7]};
				5'd8:	res <= {a[7:0], a[31:8]};
				5'd9:	res <= {a[8:0], a[31:9]};
				5'd10:	res <= {a[9:0], a[31:10]};
				5'd11:	res <= {a[10:0], a[31:11]};
				5'd12:	res <= {a[11:0], a[31:12]};
				5'd13:	res <= {a[12:0], a[31:13]};
				5'd14:	res <= {a[13:0], a[31:14]};
				5'd15:	res <= {a[14:0], a[31:15]};
				5'd16:	res <= {a[15:0], a[31:16]};
				5'd17:	res <= {a[16:0], a[31:17]};
				5'd18:	res <= {a[17:0], a[31:18]};
				5'd19:	res <= {a[18:0], a[31:19]};
				5'd20:	res <= {a[19:0], a[31:20]};
				5'd21:	res <= {a[20:0], a[31:21]};
				5'd22:	res <= {a[21:0], a[31:22]};
				5'd23:	res <= {a[22:0], a[31:23]};
				5'd24:	res <= {a[23:0], a[31:24]};
				5'd25:	res <= {a[24:0], a[31:25]};
				5'd26:	res <= {a[25:0], a[31:26]};
				5'd27:	res <= {a[26:0], a[31:27]};
				5'd28:	res <= {a[27:0], a[31:28]};
				5'd29:	res <= {a[28:0], a[31:29]};
				5'd30:	res <= {a[29:0], a[31:30]};
				5'd31:	res <= {a[30:0], a[31]};
				default: res <= a;
			endcase
		end

endmodule
